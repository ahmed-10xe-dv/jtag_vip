package jtag_seqs_pkg;
    import jtag_pkg::*;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "jtag_sequence.sv"
    // include rest of seqs as follows//
    
endpackage