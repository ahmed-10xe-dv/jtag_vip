package jtag_tests_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import jtag_pkg::*;
    import jtag_seqs_pkg::*;
    
    `include "jtag_base_test.sv"
    // include rest of tests as follows//
    
endpackage